`ifndef __PANDA_EXT_DEFINES_H
`define __PANDA_EXT_DEFINES_H

typedef enum bit[1:0]{
	INT8 = 2'b00,
	INT16 = 2'b01,
	FP16 = 2'b10
}calfmt_t;

`endif
