`ifndef __UTILS_H

`define __UTILS_H

import "DPI-C" function int unsigned encode_fp16(input real d);
import "DPI-C" function real decode_fp16(input int unsigned fp16);
	
`endif
